library verilog;
use verilog.vl_types.all;
entity quanta_vlg_vec_tst is
end quanta_vlg_vec_tst;
