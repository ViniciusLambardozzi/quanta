library verilog;
use verilog.vl_types.all;
entity quanta2_vlg_vec_tst is
end quanta2_vlg_vec_tst;
